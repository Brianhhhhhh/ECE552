module insCache(clk, rst, address, dataOut, readEn, miss);
	input clk, rst, readEn;
	input [15:0] address;
	output [15:0] dataOut;
	output miss;
	
	
	
endmodule