module ALU(out, In1, In2, );

endmodule